library ieee;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;

use work.riscy_package.all;

entity extender is
  port (
    clock
  ) ;
end extender;

architecture arch of extender is

    signal 

begin

end arch ; -- arch