../../src/de0Test.vhd